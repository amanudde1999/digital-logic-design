----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Shyama Gandhi, Amro Amanuddein and Ahmed Ahmed
-- 
-- Create Date: 10/06/2021 02:31:27 PM
-- Design Name: 
-- Module Name: full_adder_2bit - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity full_adder_1bit is
    Port ( a : in STD_LOGIC;
           b : in STD_LOGIC;
           c_in : in STD_LOGIC;
           sum : out STD_LOGIC;
           c_out : out STD_LOGIC);
end full_adder_1bit;

architecture Behavioral of full_adder_1bit is

begin

sum <= a xor b xor c_in;
c_out <= (a and b) or (b and c_in) or (c_in and a);

end Behavioral;
